package RVfmt_pkg is

	type FORMAT_RV is (R_type, I_type, S_type, SB_type, U_type, UJ_type);

end RVfmt_pkg;